// Android2FPGAMemoryMap.v

// Generated using ACDS version 12.1 177 at 2013.04.22.02:29:39

`timescale 1 ps / 1 ps
module Android2FPGAMemoryMap (
		output wire [7:0] pio_export,                                 //                                  pio.export
		input  wire       reset_reset_n,                              //                                reset.reset_n
		output wire       st_bytes_to_packets_in_bytes_stream_ready,  //  st_bytes_to_packets_in_bytes_stream.ready
		input  wire       st_bytes_to_packets_in_bytes_stream_valid,  //                                     .valid
		input  wire [7:0] st_bytes_to_packets_in_bytes_stream_data,   //                                     .data
		input  wire       clk_clk,                                    //                                  clk.clk
		input  wire       st_packets_to_bytes_out_bytes_stream_ready, // st_packets_to_bytes_out_bytes_stream.ready
		output wire       st_packets_to_bytes_out_bytes_stream_valid, //                                     .valid
		output wire [7:0] st_packets_to_bytes_out_bytes_stream_data   //                                     .data
	);

	wire         packets_to_master_out_stream_endofpacket;                                           // packets_to_master:out_endofpacket -> st_packets_to_bytes_ca:in_endofpacket
	wire         packets_to_master_out_stream_valid;                                                 // packets_to_master:out_valid -> st_packets_to_bytes_ca:in_valid
	wire         packets_to_master_out_stream_startofpacket;                                         // packets_to_master:out_startofpacket -> st_packets_to_bytes_ca:in_startofpacket
	wire   [7:0] packets_to_master_out_stream_data;                                                  // packets_to_master:out_data -> st_packets_to_bytes_ca:in_data
	wire         packets_to_master_out_stream_ready;                                                 // st_packets_to_bytes_ca:in_ready -> packets_to_master:out_ready
	wire         st_packets_to_bytes_ca_out_endofpacket;                                             // st_packets_to_bytes_ca:out_endofpacket -> st_packets_to_bytes:in_endofpacket
	wire         st_packets_to_bytes_ca_out_valid;                                                   // st_packets_to_bytes_ca:out_valid -> st_packets_to_bytes:in_valid
	wire         st_packets_to_bytes_ca_out_startofpacket;                                           // st_packets_to_bytes_ca:out_startofpacket -> st_packets_to_bytes:in_startofpacket
	wire   [7:0] st_packets_to_bytes_ca_out_data;                                                    // st_packets_to_bytes_ca:out_data -> st_packets_to_bytes:in_data
	wire   [7:0] st_packets_to_bytes_ca_out_channel;                                                 // st_packets_to_bytes_ca:out_channel -> st_packets_to_bytes:in_channel
	wire         st_packets_to_bytes_ca_out_ready;                                                   // st_packets_to_bytes:in_ready -> st_packets_to_bytes_ca:out_ready
	wire         st_bytes_to_packets_out_packets_stream_endofpacket;                                 // st_bytes_to_packets:out_endofpacket -> st_bytes_to_packets_ca:in_endofpacket
	wire         st_bytes_to_packets_out_packets_stream_valid;                                       // st_bytes_to_packets:out_valid -> st_bytes_to_packets_ca:in_valid
	wire         st_bytes_to_packets_out_packets_stream_startofpacket;                               // st_bytes_to_packets:out_startofpacket -> st_bytes_to_packets_ca:in_startofpacket
	wire   [7:0] st_bytes_to_packets_out_packets_stream_data;                                        // st_bytes_to_packets:out_data -> st_bytes_to_packets_ca:in_data
	wire         st_bytes_to_packets_out_packets_stream_ready;                                       // st_bytes_to_packets_ca:in_ready -> st_bytes_to_packets:out_ready
	wire   [7:0] st_bytes_to_packets_out_packets_stream_channel;                                     // st_bytes_to_packets:out_channel -> st_bytes_to_packets_ca:in_channel
	wire         st_bytes_to_packets_ca_out_endofpacket;                                             // st_bytes_to_packets_ca:out_endofpacket -> packets_to_master:in_endofpacket
	wire         st_bytes_to_packets_ca_out_valid;                                                   // st_bytes_to_packets_ca:out_valid -> packets_to_master:in_valid
	wire         st_bytes_to_packets_ca_out_startofpacket;                                           // st_bytes_to_packets_ca:out_startofpacket -> packets_to_master:in_startofpacket
	wire   [7:0] st_bytes_to_packets_ca_out_data;                                                    // st_bytes_to_packets_ca:out_data -> packets_to_master:in_data
	wire         st_bytes_to_packets_ca_out_ready;                                                   // packets_to_master:in_ready -> st_bytes_to_packets_ca:out_ready
	wire         packets_to_master_avalon_master_waitrequest;                                        // packets_to_master_avalon_master_translator:av_waitrequest -> packets_to_master:waitrequest
	wire  [31:0] packets_to_master_avalon_master_writedata;                                          // packets_to_master:writedata -> packets_to_master_avalon_master_translator:av_writedata
	wire  [31:0] packets_to_master_avalon_master_address;                                            // packets_to_master:address -> packets_to_master_avalon_master_translator:av_address
	wire         packets_to_master_avalon_master_write;                                              // packets_to_master:write -> packets_to_master_avalon_master_translator:av_write
	wire         packets_to_master_avalon_master_read;                                               // packets_to_master:read -> packets_to_master_avalon_master_translator:av_read
	wire  [31:0] packets_to_master_avalon_master_readdata;                                           // packets_to_master_avalon_master_translator:av_readdata -> packets_to_master:readdata
	wire   [3:0] packets_to_master_avalon_master_byteenable;                                         // packets_to_master:byteenable -> packets_to_master_avalon_master_translator:av_byteenable
	wire         packets_to_master_avalon_master_readdatavalid;                                      // packets_to_master_avalon_master_translator:av_readdatavalid -> packets_to_master:readdatavalid
	wire         packets_to_master_avalon_master_translator_avalon_universal_master_0_waitrequest;   // pio_s1_translator:uav_waitrequest -> packets_to_master_avalon_master_translator:uav_waitrequest
	wire   [2:0] packets_to_master_avalon_master_translator_avalon_universal_master_0_burstcount;    // packets_to_master_avalon_master_translator:uav_burstcount -> pio_s1_translator:uav_burstcount
	wire  [31:0] packets_to_master_avalon_master_translator_avalon_universal_master_0_writedata;     // packets_to_master_avalon_master_translator:uav_writedata -> pio_s1_translator:uav_writedata
	wire  [31:0] packets_to_master_avalon_master_translator_avalon_universal_master_0_address;       // packets_to_master_avalon_master_translator:uav_address -> pio_s1_translator:uav_address
	wire         packets_to_master_avalon_master_translator_avalon_universal_master_0_lock;          // packets_to_master_avalon_master_translator:uav_lock -> pio_s1_translator:uav_lock
	wire         packets_to_master_avalon_master_translator_avalon_universal_master_0_write;         // packets_to_master_avalon_master_translator:uav_write -> pio_s1_translator:uav_write
	wire         packets_to_master_avalon_master_translator_avalon_universal_master_0_read;          // packets_to_master_avalon_master_translator:uav_read -> pio_s1_translator:uav_read
	wire  [31:0] packets_to_master_avalon_master_translator_avalon_universal_master_0_readdata;      // pio_s1_translator:uav_readdata -> packets_to_master_avalon_master_translator:uav_readdata
	wire         packets_to_master_avalon_master_translator_avalon_universal_master_0_debugaccess;   // packets_to_master_avalon_master_translator:uav_debugaccess -> pio_s1_translator:uav_debugaccess
	wire   [3:0] packets_to_master_avalon_master_translator_avalon_universal_master_0_byteenable;    // packets_to_master_avalon_master_translator:uav_byteenable -> pio_s1_translator:uav_byteenable
	wire         packets_to_master_avalon_master_translator_avalon_universal_master_0_readdatavalid; // pio_s1_translator:uav_readdatavalid -> packets_to_master_avalon_master_translator:uav_readdatavalid
	wire  [31:0] pio_s1_translator_avalon_anti_slave_0_writedata;                                    // pio_s1_translator:av_writedata -> pio:writedata
	wire   [1:0] pio_s1_translator_avalon_anti_slave_0_address;                                      // pio_s1_translator:av_address -> pio:address
	wire         pio_s1_translator_avalon_anti_slave_0_chipselect;                                   // pio_s1_translator:av_chipselect -> pio:chipselect
	wire         pio_s1_translator_avalon_anti_slave_0_write;                                        // pio_s1_translator:av_write -> pio:write_n
	wire  [31:0] pio_s1_translator_avalon_anti_slave_0_readdata;                                     // pio:readdata -> pio_s1_translator:av_readdata
	wire         rst_controller_reset_out_reset;                                                     // rst_controller:reset_out -> [packets_to_master:reset_n, packets_to_master_avalon_master_translator:reset, pio:reset_n, pio_s1_translator:reset, st_bytes_to_packets:reset_n, st_bytes_to_packets_ca:reset_n, st_packets_to_bytes:reset_n, st_packets_to_bytes_ca:reset_n]

	altera_avalon_packets_to_master #(
		.FAST_VER    (0),
		.FIFO_DEPTHS (2),
		.FIFO_WIDTHU (1)
	) packets_to_master (
		.clk               (clk_clk),                                       //           clk.clk
		.reset_n           (~rst_controller_reset_out_reset),               //     clk_reset.reset_n
		.out_ready         (packets_to_master_out_stream_ready),            //    out_stream.ready
		.out_valid         (packets_to_master_out_stream_valid),            //              .valid
		.out_data          (packets_to_master_out_stream_data),             //              .data
		.out_startofpacket (packets_to_master_out_stream_startofpacket),    //              .startofpacket
		.out_endofpacket   (packets_to_master_out_stream_endofpacket),      //              .endofpacket
		.in_ready          (st_bytes_to_packets_ca_out_ready),              //     in_stream.ready
		.in_valid          (st_bytes_to_packets_ca_out_valid),              //              .valid
		.in_data           (st_bytes_to_packets_ca_out_data),               //              .data
		.in_startofpacket  (st_bytes_to_packets_ca_out_startofpacket),      //              .startofpacket
		.in_endofpacket    (st_bytes_to_packets_ca_out_endofpacket),        //              .endofpacket
		.address           (packets_to_master_avalon_master_address),       // avalon_master.address
		.readdata          (packets_to_master_avalon_master_readdata),      //              .readdata
		.read              (packets_to_master_avalon_master_read),          //              .read
		.write             (packets_to_master_avalon_master_write),         //              .write
		.writedata         (packets_to_master_avalon_master_writedata),     //              .writedata
		.waitrequest       (packets_to_master_avalon_master_waitrequest),   //              .waitrequest
		.readdatavalid     (packets_to_master_avalon_master_readdatavalid), //              .readdatavalid
		.byteenable        (packets_to_master_avalon_master_byteenable)     //              .byteenable
	);

	altera_avalon_st_bytes_to_packets #(
		.CHANNEL_WIDTH (8),
		.ENCODING      (0)
	) st_bytes_to_packets (
		.clk               (clk_clk),                                              //                clk.clk
		.reset_n           (~rst_controller_reset_out_reset),                      //          clk_reset.reset_n
		.out_channel       (st_bytes_to_packets_out_packets_stream_channel),       // out_packets_stream.channel
		.out_ready         (st_bytes_to_packets_out_packets_stream_ready),         //                   .ready
		.out_valid         (st_bytes_to_packets_out_packets_stream_valid),         //                   .valid
		.out_data          (st_bytes_to_packets_out_packets_stream_data),          //                   .data
		.out_startofpacket (st_bytes_to_packets_out_packets_stream_startofpacket), //                   .startofpacket
		.out_endofpacket   (st_bytes_to_packets_out_packets_stream_endofpacket),   //                   .endofpacket
		.in_ready          (st_bytes_to_packets_in_bytes_stream_ready),            //    in_bytes_stream.ready
		.in_valid          (st_bytes_to_packets_in_bytes_stream_valid),            //                   .valid
		.in_data           (st_bytes_to_packets_in_bytes_stream_data)              //                   .data
	);

	altera_avalon_st_packets_to_bytes #(
		.CHANNEL_WIDTH (8),
		.ENCODING      (0)
	) st_packets_to_bytes (
		.clk              (clk_clk),                                    //               clk.clk
		.reset_n          (~rst_controller_reset_out_reset),            //         clk_reset.reset_n
		.in_ready         (st_packets_to_bytes_ca_out_ready),           // in_packets_stream.ready
		.in_valid         (st_packets_to_bytes_ca_out_valid),           //                  .valid
		.in_data          (st_packets_to_bytes_ca_out_data),            //                  .data
		.in_channel       (st_packets_to_bytes_ca_out_channel),         //                  .channel
		.in_startofpacket (st_packets_to_bytes_ca_out_startofpacket),   //                  .startofpacket
		.in_endofpacket   (st_packets_to_bytes_ca_out_endofpacket),     //                  .endofpacket
		.out_ready        (st_packets_to_bytes_out_bytes_stream_ready), //  out_bytes_stream.ready
		.out_valid        (st_packets_to_bytes_out_bytes_stream_valid), //                  .valid
		.out_data         (st_packets_to_bytes_out_bytes_stream_data)   //                  .data
	);

	Android2FPGAMemoryMap_pio pio (
		.clk        (clk_clk),                                          //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                  //               reset.reset_n
		.address    (pio_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~pio_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (pio_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (pio_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (pio_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.out_port   (pio_export)                                        // external_connection.export
	);

	Android2FPGAMemoryMap_st_packets_to_bytes_ca st_packets_to_bytes_ca (
		.clk               (clk_clk),                                    //   clk.clk
		.reset_n           (~rst_controller_reset_out_reset),            // reset.reset_n
		.in_ready          (packets_to_master_out_stream_ready),         //    in.ready
		.in_valid          (packets_to_master_out_stream_valid),         //      .valid
		.in_data           (packets_to_master_out_stream_data),          //      .data
		.in_startofpacket  (packets_to_master_out_stream_startofpacket), //      .startofpacket
		.in_endofpacket    (packets_to_master_out_stream_endofpacket),   //      .endofpacket
		.out_ready         (st_packets_to_bytes_ca_out_ready),           //   out.ready
		.out_valid         (st_packets_to_bytes_ca_out_valid),           //      .valid
		.out_data          (st_packets_to_bytes_ca_out_data),            //      .data
		.out_startofpacket (st_packets_to_bytes_ca_out_startofpacket),   //      .startofpacket
		.out_endofpacket   (st_packets_to_bytes_ca_out_endofpacket),     //      .endofpacket
		.out_channel       (st_packets_to_bytes_ca_out_channel)          //      .channel
	);

	Android2FPGAMemoryMap_st_bytes_to_packets_ca st_bytes_to_packets_ca (
		.clk               (clk_clk),                                              //   clk.clk
		.reset_n           (~rst_controller_reset_out_reset),                      // reset.reset_n
		.in_ready          (st_bytes_to_packets_out_packets_stream_ready),         //    in.ready
		.in_valid          (st_bytes_to_packets_out_packets_stream_valid),         //      .valid
		.in_data           (st_bytes_to_packets_out_packets_stream_data),          //      .data
		.in_channel        (st_bytes_to_packets_out_packets_stream_channel),       //      .channel
		.in_startofpacket  (st_bytes_to_packets_out_packets_stream_startofpacket), //      .startofpacket
		.in_endofpacket    (st_bytes_to_packets_out_packets_stream_endofpacket),   //      .endofpacket
		.out_ready         (st_bytes_to_packets_ca_out_ready),                     //   out.ready
		.out_valid         (st_bytes_to_packets_ca_out_valid),                     //      .valid
		.out_data          (st_bytes_to_packets_ca_out_data),                      //      .data
		.out_startofpacket (st_bytes_to_packets_ca_out_startofpacket),             //      .startofpacket
		.out_endofpacket   (st_bytes_to_packets_ca_out_endofpacket)                //      .endofpacket
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (32),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (32),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (1),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (1),
		.USE_WAITREQUEST             (1),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) packets_to_master_avalon_master_translator (
		.clk                   (clk_clk),                                                                            //                       clk.clk
		.reset                 (rst_controller_reset_out_reset),                                                     //                     reset.reset
		.uav_address           (packets_to_master_avalon_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount        (packets_to_master_avalon_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read              (packets_to_master_avalon_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write             (packets_to_master_avalon_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest       (packets_to_master_avalon_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid     (packets_to_master_avalon_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable        (packets_to_master_avalon_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata          (packets_to_master_avalon_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata         (packets_to_master_avalon_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock              (packets_to_master_avalon_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess       (packets_to_master_avalon_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address            (packets_to_master_avalon_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest        (packets_to_master_avalon_master_waitrequest),                                        //                          .waitrequest
		.av_byteenable         (packets_to_master_avalon_master_byteenable),                                         //                          .byteenable
		.av_read               (packets_to_master_avalon_master_read),                                               //                          .read
		.av_readdata           (packets_to_master_avalon_master_readdata),                                           //                          .readdata
		.av_readdatavalid      (packets_to_master_avalon_master_readdatavalid),                                      //                          .readdatavalid
		.av_write              (packets_to_master_avalon_master_write),                                              //                          .write
		.av_writedata          (packets_to_master_avalon_master_writedata),                                          //                          .writedata
		.av_burstcount         (1'b1),                                                                               //               (terminated)
		.av_beginbursttransfer (1'b0),                                                                               //               (terminated)
		.av_begintransfer      (1'b0),                                                                               //               (terminated)
		.av_chipselect         (1'b0),                                                                               //               (terminated)
		.av_lock               (1'b0),                                                                               //               (terminated)
		.av_debugaccess        (1'b0),                                                                               //               (terminated)
		.uav_clken             (),                                                                                   //               (terminated)
		.av_clken              (1'b1)                                                                                //               (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) pio_s1_translator (
		.clk                   (clk_clk),                                                                            //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                                     //                    reset.reset
		.uav_address           (packets_to_master_avalon_master_translator_avalon_universal_master_0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (packets_to_master_avalon_master_translator_avalon_universal_master_0_burstcount),    //                         .burstcount
		.uav_read              (packets_to_master_avalon_master_translator_avalon_universal_master_0_read),          //                         .read
		.uav_write             (packets_to_master_avalon_master_translator_avalon_universal_master_0_write),         //                         .write
		.uav_waitrequest       (packets_to_master_avalon_master_translator_avalon_universal_master_0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (packets_to_master_avalon_master_translator_avalon_universal_master_0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (packets_to_master_avalon_master_translator_avalon_universal_master_0_byteenable),    //                         .byteenable
		.uav_readdata          (packets_to_master_avalon_master_translator_avalon_universal_master_0_readdata),      //                         .readdata
		.uav_writedata         (packets_to_master_avalon_master_translator_avalon_universal_master_0_writedata),     //                         .writedata
		.uav_lock              (packets_to_master_avalon_master_translator_avalon_universal_master_0_lock),          //                         .lock
		.uav_debugaccess       (packets_to_master_avalon_master_translator_avalon_universal_master_0_debugaccess),   //                         .debugaccess
		.av_address            (pio_s1_translator_avalon_anti_slave_0_address),                                      //      avalon_anti_slave_0.address
		.av_write              (pio_s1_translator_avalon_anti_slave_0_write),                                        //                         .write
		.av_readdata           (pio_s1_translator_avalon_anti_slave_0_readdata),                                     //                         .readdata
		.av_writedata          (pio_s1_translator_avalon_anti_slave_0_writedata),                                    //                         .writedata
		.av_chipselect         (pio_s1_translator_avalon_anti_slave_0_chipselect),                                   //                         .chipselect
		.av_read               (),                                                                                   //              (terminated)
		.av_begintransfer      (),                                                                                   //              (terminated)
		.av_beginbursttransfer (),                                                                                   //              (terminated)
		.av_burstcount         (),                                                                                   //              (terminated)
		.av_byteenable         (),                                                                                   //              (terminated)
		.av_readdatavalid      (1'b0),                                                                               //              (terminated)
		.av_waitrequest        (1'b0),                                                                               //              (terminated)
		.av_writebyteenable    (),                                                                                   //              (terminated)
		.av_lock               (),                                                                                   //              (terminated)
		.av_clken              (),                                                                                   //              (terminated)
		.uav_clken             (1'b0),                                                                               //              (terminated)
		.av_debugaccess        (),                                                                                   //              (terminated)
		.av_outputenable       ()                                                                                    //              (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (1),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2)
	) rst_controller (
		.reset_in0  (~reset_reset_n),                 // reset_in0.reset
		.clk        (clk_clk),                        //       clk.clk
		.reset_out  (rst_controller_reset_out_reset), // reset_out.reset
		.reset_in1  (1'b0),                           // (terminated)
		.reset_in2  (1'b0),                           // (terminated)
		.reset_in3  (1'b0),                           // (terminated)
		.reset_in4  (1'b0),                           // (terminated)
		.reset_in5  (1'b0),                           // (terminated)
		.reset_in6  (1'b0),                           // (terminated)
		.reset_in7  (1'b0),                           // (terminated)
		.reset_in8  (1'b0),                           // (terminated)
		.reset_in9  (1'b0),                           // (terminated)
		.reset_in10 (1'b0),                           // (terminated)
		.reset_in11 (1'b0),                           // (terminated)
		.reset_in12 (1'b0),                           // (terminated)
		.reset_in13 (1'b0),                           // (terminated)
		.reset_in14 (1'b0),                           // (terminated)
		.reset_in15 (1'b0)                            // (terminated)
	);

endmodule
